module andt(
  input [7:0] a,b,
  output [7:0] y
);
  
  assign y = a & b ;
  
endmodule
